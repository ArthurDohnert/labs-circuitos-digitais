library verilog;
use verilog.vl_types.all;
entity DECOD416_vlg_vec_tst is
end DECOD416_vlg_vec_tst;
