library verilog;
use verilog.vl_types.all;
entity RCA16_vlg_vec_tst is
end RCA16_vlg_vec_tst;
