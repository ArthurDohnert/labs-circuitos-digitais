library verilog;
use verilog.vl_types.all;
entity lab07 is
    port(
        Q               : out    vl_logic;
        D               : in     vl_logic;
        clk             : in     vl_logic
    );
end lab07;
