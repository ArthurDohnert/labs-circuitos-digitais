library verilog;
use verilog.vl_types.all;
entity FSM_elevador_vlg_vec_tst is
end FSM_elevador_vlg_vec_tst;
