library verilog;
use verilog.vl_types.all;
entity CodificadordePrioridade_vlg_vec_tst is
end CodificadordePrioridade_vlg_vec_tst;
