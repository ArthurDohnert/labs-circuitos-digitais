library verilog;
use verilog.vl_types.all;
entity lab07_vlg_vec_tst is
end lab07_vlg_vec_tst;
