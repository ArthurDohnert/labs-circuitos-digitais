library verilog;
use verilog.vl_types.all;
entity RCA4_vlg_vec_tst is
end RCA4_vlg_vec_tst;
