library verilog;
use verilog.vl_types.all;
entity UnidadeAritmetica_vlg_vec_tst is
end UnidadeAritmetica_vlg_vec_tst;
